interface FFT4If;    
    logic [15:0] x0_re, x0_im, x1_re, x1_im, x2_re, x2_im, x3_re, x3_im;
    logic [15:0] y0_re, y0_im, y1_re, y1_im, y2_re, y2_im, y3_re, y3_im;
    logic clk; // Clock signal
endinterface 
